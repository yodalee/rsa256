package RSA_pkg;

parameter MOD_WIDTH = 256;

typedef logic [MOD_WIDTH-1:0] KeyType;

endpackage