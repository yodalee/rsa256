module dummy (
  input clk
);
endmodule